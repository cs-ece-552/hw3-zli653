/*
    CS/ECE 552 Spring '19
    Homework #3, Problem 2
    
    a 1-bit full adder
*/
module fullAdder_1b(A, B, C_in, S, C_out);
    input  A, B;
	input  C_in;
    output S;
    output C_out;

	// YOUR CODE HERE

endmodule
