/*
    CS/ECE 552 Spring '19
    Homework #3, Problem 1

    2-1 mux template
*/
module mux2_1(InA, InB, InC, InD, S, Out);
    input   InA, InB, InC, InD;
    input   S;
    output  Out;

    // YOUR CODE HERE

endmodule
